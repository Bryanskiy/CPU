module execute(
    input logic[(`WORD - 1):0] rdata1E, rdata2E, immE, pcE,
    input logic regWriteE, memWriteE, mem2regE,

    output logic[(`WORD - 1):0] writeDataM, writeRegM, ALUOutM,
    output logic ZeroM
);

    

endmodule