module top(
    input logic clk
);
endmodule