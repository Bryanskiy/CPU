module hazard(
    /* for bypass */
    input logic[(`REG_SIZE - 1):0] writeRegM, writeRegW,
    input logic regWriteM, regWriteW
);
endmodule