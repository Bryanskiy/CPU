module datapath();
    // next PC logic

    // register file logic

    // ALU logic
endmodule