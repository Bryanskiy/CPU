module datapath(
    input logic clk,
    input logic regWrite,
    input logic memWrite,
    input logic[3:0] ALUControl
);
    // next PC logic

    // register file logic

    // ALU logic
endmodule